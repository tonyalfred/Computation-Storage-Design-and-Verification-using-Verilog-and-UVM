/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         comp_strg_defines.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

  `ifndef COMP_STRG_DEFINES
    `define COMP_STRG_DEFINES

    `ifndef STRG_DATA_WIDTH
      `define STRG_DATA_WIDTH     32
    `endif

    `ifndef STRG_ADDRESS_WIDTH
      `define STRG_ADDRESS_WIDTH  10
    `endif 
  `endif

/**********************************************************************************************************************
*  END OF FILE: comp_strg_defines.sv
*********************************************************************************************************************/