/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         comp_strg_types.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

`ifndef COMP_STRG_TYPES
  `define COMP_STRG_TYPES
    
  typedef enum bit [2:0] {READ = 0, WRITE = 1, ADD = 2, SUB = 3, NOP = 4} comp_strg_transaction_type_t;

`endif

/**********************************************************************************************************************
*  END OF FILE: comp_strg_types.sv
*********************************************************************************************************************/